
module PreLab_3_2BitAdder_tb();

//inputs into PreLab tests
reg x_0, x_1, y_0, y_1;

wire S, C_1, C_2;

PreLab_3_2BitAdder tg1(.x_0(x_0), .x_1(x_1), .y_0(y_0), .y_1(y_1), .S(S), .C_1(C_1), .C_2(C_2) );

initial begin

  x_1 = 0; x_0 = 0; y_1 = 0; y_0 = 0; #100;

  x_1 = 0; x_0 = 0; y_1 = 0; y_0 = 1; #100;

  x_1 = 0; x_0 = 0; y_1 = 1; y_0 = 0; #100;

  x_1 = 0; x_0 = 0; y_1 = 1; y_0 = 1; #100;

  x_1 = 0; x_0 = 1; y_1 = 0; y_0 = 0; #100;

  x_1 = 0; x_0 = 1; y_1 = 0; y_0 = 1; #100;

  x_1 = 0; x_0 = 1; y_1 = 1; y_0 = 0; #100;

  x_1 = 0; x_0 = 1; y_1 = 1; y_0 = 1; #100;

  x_1 = 1; x_0 = 0; y_1 = 0; y_0 = 0; #100;

  x_1 = 1; x_0 = 0; y_1 = 0; y_0 = 1; #100;

  x_1 = 1; x_0 = 0; y_1 = 1; y_0 = 0; #100;

  x_1 = 1; x_0 = 0; y_1 = 1; y_0 = 1; #100;

  x_1 = 1; x_0 = 1; y_1 = 0; y_0 = 0; #100;

  x_1 = 1; x_0 = 1; y_1 = 0; y_0 = 1; #100;

  x_1 = 1; x_0 = 1; y_1 = 1; y_0 = 0; #100;

  x_1 = 1; x_0 = 1; y_1 = 1; y_0 = 1; #100;

end

endmodule
